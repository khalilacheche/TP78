architecture rtl of led_driver is
    --ok: "000000000000" &
    --    "000000000000" &
    --    "000001010100" &
    --    "000010110100" &
    --    "000010111000" &
    --    "000010110100" &
    --    "000001010100" &
    --    "000000000000" &
    --    "000000000000";
begin
end architecture rtl;
