architecture rtl of debouncer is
begin
end architecture rtl; 
