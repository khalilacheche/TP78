architecture rtl of led_driver is
  constant ok : std_logic_vector(107 downto 0):=
     "000000000000" &
     "000000000000" &
     "000001010100" &
     "000010110100" &
     "000010111000" &
     "000010110100" &
     "000001010100" &
     "000000000000" &
     "000000000000";

    constant fr : std_logic_vector(107 downto 0):=
        "000000000000" &
        "000000000000" &
        "000011100000" &
        "000010010000" &
        "000011011000" &
        "000010010000" &
        "000010010100" &
        "000000000000" &
        "000000000000";

    constant cup : std_logic_vector(107 downto 0):=
        "000000000000" &
        "000000000000" &
        "000000000000" &
        "000011000111" &
        "000010101101" &
        "000010101111" &
        "000011111100" &
        "000000000100" &
        "000000000000";
    constant drink : std_logic_vector(107 downto 0):=
        "000000000000" &
        "000000000000" &
        "001000000000" &
        "001101000100" &
        "111110111101" &
        "101101101110" &
        "111101101101" &
        "000000000000" &
        "000000000000";
    constant x_new : std_logic_vector(107 downto 0):=
        "100000011100" &
        "000100010100" &
        "000000011100" &
        "010000010000" &
        "001000011100" &
        "010000000000" &
        "001001110101" &
        "100001010111" &
        "000101010111";
    constant donate : std_logic_vector(107 downto 0):=
        "001011100000" &
        "010110100000" &
        "010110111100" &
        "010100001010" &
        "001001111101" &
        "001000111111" &
        "111001011100" &
        "101001111011" &
        "111000000000";
begin
  process(msg, progress_led)
    begin
    case msg is
    when "001" =>
    leds <= fr; --fr
    when "010" =>
    leds <= drink; --drink
    when "011" =>
    leds <= x_new; --x_new
    when "100" =>
    leds <= cup; --cup
    when "101" =>
    leds <= donate; --donate
    when "110" =>
      leds<= ok;
      case(change_count_2) is
        when "00001" => leds(11)<='1';
        when "00010" => leds(11)<='1'; leds(11+1*12)<='1';
        when "00011" =>leds(11)<='1'; leds(11+1*12)<='1'; leds(11+2*12)<='1';
        when "00100" =>leds(11)<='1'; leds(11+1*12)<='1';leds(11+2*12)<='1'; leds(11+3*12)<='1';
        when "00101" =>leds(11)<='1';leds(11+1*12)<='1';leds(11+2*12)<='1';leds(11+3*12)<='1';leds(11+4*12)<='1';
        when "00110" =>leds(11)<='1';leds(11+1*12)<='1';leds(11+2*12)<='1';leds(11+3*12)<='1';leds(11+4*12)<='1';leds(11+5*12)<='1';
        when "00111" =>leds(11)<='1';leds(11+1*12)<='1';leds(11+2*12)<='1';leds(11+3*12)<='1';leds(11+4*12)<='1';leds(11+5*12)<='1';leds(11+6*12)<='1';
        when "01000" =>leds(11)<='1';leds(11+1*12)<='1';leds(11+2*12)<='1';leds(11+3*12)<='1';leds(11+4*12)<='1';leds(11+5*12)<='1';leds(11+6*12)<='1';leds(11+7*12)<='1';
        when "01001" =>leds(11)<='1';leds(11+1*12)<='1';leds(11+2*12)<='1';leds(11+3*12)<='1';leds(11+4*12)<='1';leds(11+5*12)<='1';leds(11+6*12)<='1';leds(11+7*12)<='1'; leds(11+8*12)<='1';
        when others =>
      end case;
      case(change_count_1) is
        when "00001" => leds(10)<='1';
        when "00010" => leds(10)<='1'; leds(10+1*12)<='1';
        when "00011" =>leds(10)<='1'; leds(10+1*12)<='1'; leds(10+2*12)<='1';
        when "00100" =>leds(10)<='1'; leds(10+1*12)<='1';leds(10+2*12)<='1'; leds(10+3*12)<='1';
        when "00101" =>leds(10)<='1';leds(10+1*12)<='1';leds(10+2*12)<='1';leds(10+3*12)<='1';leds(10+4*12)<='1';
        when "00110" =>leds(10)<='1';leds(10+1*12)<='1';leds(10+2*12)<='1';leds(10+3*12)<='1';leds(10+4*12)<='1';leds(10+5*12)<='1';
        when "00111" =>leds(10)<='1';leds(10+1*12)<='1';leds(10+2*12)<='1';leds(10+3*12)<='1';leds(10+4*12)<='1';leds(10+5*12)<='1';leds(10+6*12)<='1';
        when "01000" =>leds(10)<='1';leds(10+1*12)<='1';leds(10+2*12)<='1';leds(10+3*12)<='1';leds(10+4*12)<='1';leds(10+5*12)<='1';leds(10+6*12)<='1';leds(10+7*12)<='1';
        when "01001" =>leds(10)<='1';leds(10+1*12)<='1';leds(10+2*12)<='1';leds(10+3*12)<='1';leds(10+4*12)<='1';leds(10+5*12)<='1';leds(10+6*12)<='1';leds(10+7*12)<='1'; leds(10+8*12)<='1';
        when others =>
      end case;
      case(change_count_05) is
        when "00001" => leds(9)<='1';
        when "00010" => leds(9)<='1'; leds(9+1*12)<='1';
        when "00011" =>leds(9)<='1'; leds(9+1*12)<='1'; leds(9+2*12)<='1';
        when "00100" =>leds(9)<='1'; leds(9+1*12)<='1';leds(9+2*12)<='1'; leds(9+3*12)<='1';
        when "00101" =>leds(9)<='1';leds(9+1*12)<='1';leds(9+2*12)<='1';leds(9+3*12)<='1';leds(9+4*12)<='1';
        when "00110" =>leds(9)<='1';leds(9+1*12)<='1';leds(9+2*12)<='1';leds(9+3*12)<='1';leds(9+4*12)<='1';leds(9+5*12)<='1';
        when "00111" =>leds(9)<='1';leds(9+1*12)<='1';leds(9+2*12)<='1';leds(9+3*12)<='1';leds(9+4*12)<='1';leds(9+5*12)<='1';leds(9+6*12)<='1';
        when "01000" =>leds(9)<='1';leds(9+1*12)<='1';leds(9+2*12)<='1';leds(9+3*12)<='1';leds(9+4*12)<='1';leds(9+5*12)<='1';leds(9+6*12)<='1';leds(9+7*12)<='1';
        when "01001" =>leds(9)<='1';leds(9+1*12)<='1';leds(9+2*12)<='1';leds(9+3*12)<='1';leds(9+4*12)<='1';leds(9+5*12)<='1';leds(9+6*12)<='1';leds(9+7*12)<='1'; leds(9+8*12)<='1';
        when others =>
      end case;
      case(change_count_02) is
        when "00001" => leds(8)<='1';
        when "00010" => leds(8)<='1'; leds(8+1*12)<='1';
        when "00011" =>leds(8)<='1'; leds(8+1*12)<='1'; leds(8+2*12)<='1';
        when "00100" =>leds(8)<='1'; leds(8+1*12)<='1';leds(8+2*12)<='1'; leds(8+3*12)<='1';
        when "00101" =>leds(8)<='1';leds(8+1*12)<='1';leds(8+2*12)<='1';leds(8+3*12)<='1';leds(8+4*12)<='1';
        when "00110" =>leds(8)<='1';leds(8+1*12)<='1';leds(8+2*12)<='1';leds(8+3*12)<='1';leds(8+4*12)<='1';leds(8+5*12)<='1';
        when "00111" =>leds(8)<='1';leds(8+1*12)<='1';leds(8+2*12)<='1';leds(8+3*12)<='1';leds(8+4*12)<='1';leds(8+5*12)<='1';leds(8+6*12)<='1';
        when "01000" =>leds(8)<='1';leds(8+1*12)<='1';leds(8+2*12)<='1';leds(8+3*12)<='1';leds(8+4*12)<='1';leds(8+5*12)<='1';leds(8+6*12)<='1';leds(8+7*12)<='1';
        when "01001" =>leds(8)<='1';leds(8+1*12)<='1';leds(8+2*12)<='1';leds(8+3*12)<='1';leds(8+4*12)<='1';leds(8+5*12)<='1';leds(8+6*12)<='1';leds(8+7*12)<='1'; leds(8+8*12)<='1';
        when others =>
      end case;
    --leds <= ok + change
    when "111" =>
    leds(0)<= progress_led;
    leds(107 downto 1)<= std_logic_vector(to_unsigned(0,107));
    when others =>
    leds <= std_logic_vector(to_unsigned(0,108)); --off
    end case;
end process;
end architecture rtl;
