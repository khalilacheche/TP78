architecture rtl of drink_preparation is
--Preparation times are as follows (ordered from MSB to LSB):
--5, 7, 7, 9, 13
--Prices are as follows (ordered from MSB to LSB):
--1.2, 1.4, 1.4, 1.8, 2.5
--You may use the >>float_to_fixed<< routine to convert to unsigned.
--Numbers of ingredients packages are as follows (ordered from MSB to LSB):
--2, 2, 2, 2, 1
begin
end architecture rtl;
