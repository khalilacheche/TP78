architecture rtl of storage_ctl is
begin
end architecture rtl;
