architecture rtl of timed_button is
begin
end architecture rtl;
