architecture rtl of money_storage is
begin
end architecture rtl; 
