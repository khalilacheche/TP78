architecture rtl of main_fsm is
begin
end architecture rtl;
