architecture rtl of disp_driver is
begin
end architecture rtl;
