architecture rtl of machine is
begin
end architecture rtl;
