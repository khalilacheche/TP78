architecture rtl of timer is
begin
end architecture rtl;
