architecture rtl of sum_splitter is
begin
end architecture rtl;
