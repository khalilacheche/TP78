architecture rtl of bin_to_bcd is
    --It is guaranteed that bin never exceeds two digits, i.e., 99.
begin
end architecture rtl;
